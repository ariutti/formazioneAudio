BZh91AY&SYR�+% ߀Px��g߰����P�z�v1�a$I���dd'��Ҟ���d ���"!<���2h���2d0 4" � 6@�� �4���L� �LL&4��%552���=�OH =@A�%c�I��W�a"��3
��.��6�ؿ	@,M ������Wd��p���:4O�����2�ߏEb�>vG�]�lۙ%`�l#OU�Fi�)�jJơc
�$�T
�!�4��,�	óZK-R\�PxN]FE8!(���K��ic��N�q���sܮ:�b��&�vO��xi��.#�6�����m��3_B�r�k��5�ʕR�Yc|̍.��\	!2����b�GL�Q���>'f��ޘ���*�m� ��n�d������C\��5< G4�.�Q������P�0�Ҳ��m���d��v�ԑ �zd��[6�=VXU����K�c<�:(��;���؈ߴ���Gv[���w^mst)���.�p�Q8�L0������c� ����Ar���#���9�6.,���!���<sLTLV�n*Y�B�*3��1�����G�~�S��L�|Ӆq���Ԙ�sQ����H#)Hi鼵j&Z��$^n�g=Y�r��2oeD%q��	���{��Z���qI���t3��ܮPA��ĥ��JD=�D2 �<!�­�er�X��j@�xM��hQ�U�s*ʥ:!\&7��\����d=Dt�����\~��N`��j�+Res�G1f�M4F[��Z�D�&d����@��k��W
��&Q�a�*1R��]C��k�k�^ԋ�䙐tU��`�%YuZS��t�왆P�ɠ�с(L8hdz
b+�kօ�u�¨1�*#�.�dl���v}7!��딹�d�Jp���"�(H)I��