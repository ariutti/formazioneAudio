BZh91AY&SY��?�  �߀@x��g߰����P8�se�sp�)���؁F�� 4�h��b ���bh0 �i�10��B4�@���M hH�L`�a4� d�@�I��#ڈ����=SOP=@d4 h��$4
�B߰��e0lI���$]�jj�+5v��J��$nÂ��.�/2>��ƞv@NEk������c����%�9�/u�Yi�����{�೰�S�y�l;zIF�p�q���4�k����]|5��Fj�U��mm����7��Ey��O���;�MF4y�&�9�,�w+d�$��Y	�j�di��6b��	�u�{�}y/~
��%i���գ�[��Q��:�/O��Ѣx��,��0�%�D�d+	<�-��qw�����N"U&�H1*jo�_�(����H�oD"5r��Z��`����X$q�n��_;���$os����o�1�pX<Hd�q����Q��3b4�g_	�p&�G1�Q	��.������,���m`��eGw��$�U� ��$ȐᰉRD�=.��K�.:�^~ԋ�rI�8��rE�a,U�V	��E+y�/� 훈��Ã��f�A� �cH1�6�0>64J_�Ǩ��<���̌FR��9S#U-y
�c"Ó��p��}�Hn�-(�ʦ��jC98ٻ1����&e����zXaD���P�A��G�%�08��('���Nj������Ś�f����`���[$"SX�>�4UbJ��)�
ӎ(֌��"Zg+���L��T�i���a-d+�ز{�
���R}*񍁠��7���"�(H{J�� 