BZh91AY&SY�'	r  �߀Px��g߰����P>���vͰI�F�AM���Fj4�C& IM54jjoJ�=F�    �D�S�M2z��    9�L�����a0CLM0D�eM��j��@  �h  �\$:��N���}�S0&df���yii�������c��k��8�3��B����f����!��b���D� P��J�p�N����j��CV�\�N�)���	$ Y��g 6�����ai�,qc�VPy����h�W(��jވW�	c�I$ G�Ax�,XjeR�g1"��1���)$*wz)5�v�B�c�"�E�:��V���D�Vv~�c=ͼ�� GD�<��g�L�ܚ�k�1lڌ�a�e;	���Y�����P�T��k�nuk��1����1ft��M�&��Ck�gJi\�ut%�Po�F��B���O�������8<c���T�A�@�`C�QaS.����&��R�$�j�r��]E���X�!�_<�ws�d�:_�3T#�%z��bќ�Yo.$�8	-�+�nً�OI&ꨅne����ĵl=��p��biZ��Q����H����0�g�H'q�@��%���Gl�2-t�D��ZɆ�uZ�g5U�=� ��Cs>�	ud&ȶ1���P|pO�K�Rr�v��6���7#�^^�P��׼1 @��4g����j�����2ةD1_� A�R��L�.��t[����J����,��u�X�^W�U�����f&P�&6U}�+>R0�!��Y���tkfE�3�GcHa����
?��H�
��.@