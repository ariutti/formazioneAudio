BZh91AY&SY�$ _�Px��g߰?���P�r�q�i���ҙ���4�Q��M4f�� 4�MH4��A�     !!ML��'��&�  �0��	��i� ɦ���C$�&C=��4�@6�P��$B
��/x��u����d��6/�rP%��8?�Ԙjl���-xp9��S��E�է�J��z�?l-��cf���K,cD�ىAk�5�^x�*	%]P@\���x�wU�8�Ql2T��3S(�8b�j�y׶�_�����"�rU�2v5�C�Z�kě����y0A F�=$_cm�g^���`Η�6�O
�V�F7����;.L��
XȀv3>�*���ř�{�K��#��mP�I_��{R��:o������:GtN�o��R,�����*�k�Zq(�m[���?�M-�b��V"�brLg)�tkZǚ��|��fK�f��^<$x�{!J҈�P�V R��l����{m�
����q�[�gu���G��f��,r�D�ji։�*��_�an"��*�#�čD���#R�%pOF�ۉ�q(��#ߏ$�����,�T]j��'�3VTV�T"��o�#�a�6�DM��n�SP.O�2�Tm�$ִ���,�0o\e#�+]�il8/��	��gT�n�"2B�h�L�؆�HYm�o�F2�M���w��%H�C�^+[\[2V��1��Y���7�$"��R�����B���e��*S3�n�k����厩�R%�9�UXd;�n�)�@�Z����%D�� g-�ü���#,�=$���W �������E�R�4F� &�.XPrR��O�� 6��W��p���g��[���l+>�Cc焹��YrS���"�(H� 